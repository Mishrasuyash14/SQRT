module tbench();

wire [31:0]out;
reg [31:0]ia,ib;
new_div dut(out,ia,ib);
initial
 begin
 
 ia=0;ib=32'b00000000000000000000000000001010;
 #10 ia=32'b01000010110100100000000000000000; ib=32'b01000010010101000000000000000000;
 #10 ia=32'b01000011010101100000000000000000; ib=32'b01000010010101000000000000000000;
 #10 ia=32'b01000001110010000000000000000000; ib=32'b01000010010010000000000000000000;
 #50 $stop;
 end
endmodule
